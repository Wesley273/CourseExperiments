CIRCUIT EXP5_7
VI 1 0 AC 1V
R1 1 2 10K
R2 2 4 10K
R3 3 0 5K
C1 1 3 100PF
C2 3 4 100PF
C3 2 0 200PF
.AC LIN 100000 1MHZ 1MEGHZ
.PROBE
.END