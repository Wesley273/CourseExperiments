CIRCUIT EXP4_6
VS 1 0 DC 84V
R1 1 2 RMOD 2K
R2 2 0 RMOD 10K
G1 2 0 POLY(1) 2 0 0 0.3 0.04 0 2
.MODEL RMOD RES(R=1 TCE=0)
.TRAN 10U 4M
.PROBE
.END