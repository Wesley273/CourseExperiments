CIRCUIT EXP3_2
*VIM 3 0 SIN(10MV 50MV 500HZ 0.3MS 1E3 30DEG)
VIM 3 0 SFFM (5MV 30MV 500HZ 6 50HZ)
V1 6 0 DC 20V
R1 3 1 RMOD 50
R2 5 6 RMOD 3.5K
R3 2 0 RMOD 500K
R4 4 0 RMOD 1.5K
R5 7 0 RMOD 20K
C1 1 2 CMOD 1UF
C2 4 0 CMOD 10UF
C3 5 7 CMOD 1UF
J1 5 2 4 JNJF
.MODEL RMOD RES(R=1 TCE=0)
.MODEL LMOD IND(L=1 IL1=0 IL2=0 TC1=0 TC2=0)
.MODEL CMOD CAP(C=1 VC1=0 VC2=0 TC1=0 TC2=0)
.MODEL JNJF NJF(IS=100E-14 RD=10 RS=10 BETA=1E-3 CGD=5PF CGS=1PF VTO=-5) 
.TRAN 1US 5MS
.PROBE
.END