LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ADDER8_B IS
    PORT (
        CIN : IN STD_LOGIC;
        A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        SUM : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        COUT : OUT STD_LOGIC);
END ENTITY ADDER8_B;

ARCHITECTURE BHV OF ADDER8_B IS
    COMPONENT ADDER4 IS
        PORT (
            CIN : IN STD_LOGIC;
            A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            SUM : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            COUT : OUT STD_LOGIC);
    END COMPONENT ADDER4;
    SIGNAL DATA : STD_LOGIC_VECTOR(8 DOWNTO 0);
    SIGNAL C : STD_LOGIC;
BEGIN
    LOW : ADDER4 PORT MAP(CIN => CIN, A => A(3 DOWNTO 0), B => B(3 DOWNTO 0), COUT => C, SUM => SUM(3 DOWNTO 0));
    HIGH : ADDER4 PORT MAP(CIN => C, A => A(7 DOWNTO 4), B => B(7 DOWNTO 4), COUT => COUT, SUM => SUM(7 DOWNTO 4));
END ARCHITECTURE BHV;