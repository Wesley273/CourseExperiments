CIRCUIT EXP3_5
VI1 1 0 AC 0.5V 0DEG
VI2 2 0 AC -0.5V DEG
VDD 6 0 DC 12V
VSS 0 8 DC 12V
R1 7 0 RMOD 100K
M1 4 1 3 3 MNMOS W=20U L=5U AD=200P AS=200P
M2 5 2 3 3 MNMOS W=20U L=5U AD=200P AS=200P
M3 4 4 6 6 MPMOS W=60U L=5U AD=600P AS=600P
M4 5 4 6 6 MPMOS W=60U L=5U AD=600P AS=600P
M5 3 7 8 8 MNMOS W=20U L=5U AD=200P AS=200P
M6 7 7 8 8 MNMOS W=20U L=5U AD=200P AS=200P
.MODEL RMOD RES(R=1 TCE=0)
.MODEL LMOD IND(L=1 IL1=0 IL2=0 TC1=0 TC2=0)
.MODEL CMOD CAP(C=1 VC1=0 VC2=0 TC1=0 TC2=0)
.MODEL MNMOS NMOS(VTO=0.8 GAMMA=0.2 PHI=0.6 LAMBDA=0.03 JS=0.16 PB=0.82 CGSO=2.9E-10 CGDO=2.9E-10 CGBO=2.2E-9 RSH=6 TOX=9.5E-8 NSUB=2.5E14 XJ=1.2U LD=0.8U UO=700)
.MODEL MPMOS PMOS(VTO=-4 GAMMA=0.2 PHI=0.6 LAMBDA=0.03 JS=0.16 PB=0.82 CGSO=2.9E-10 CGDO=2.9E-10 CGBO=2.2E-9 RSH=30 TOX=9.5E-8 NSUB=1.2E14 XJ=1.0U LD=0.8U UO=235)
.AC DEC 10 1K 100MEG
.PROBE
.END