CIRCUIT EXP4_8
VIN1 1 0 DC 0V
VIN2 2 0 DC 0V
VCC1 4 0 DC 5V
VCC2 10 0 DC 5V
R1 3 4 RMOD 10K
R2 6 4 RMOD 1K
R3 4 8 RMOD 10K
R5 10 11 1K
R6 10 9 10K
Q1 5 3 1 QNPN
Q2 6 5 0 QNPN
Q3 6 7 0 QNPN
Q4 7 8 2 QNPN
Q5 12 9 6 QNPN
Q6 11 12 0 QNPN
.MODEL RMOD RES(R=1 TCE=0)
.MODEL QNPN NPN(IS=3.06E-14, BF=220 RB=0.13 RC=0.12 VAF=104 CJC=9.12P TF=0.325NS)
.TRAN 20U 2M
.PROBE
.END