LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DETECTBUCKCODE IS
    PORT (
        CLK : IN STD_LOGIC;
        BUCKIN : IN STD_LOGIC;
        RESULT : OUT STD_LOGIC
    );
END DETECTBUCKCODE;
ARCHITECTURE BHV OF DETECTBUCKCODE IS
    TYPE STATES IS(ST0, ST1, ST2, ST3, ST4, ST5, ST6);
    SIGNAL CURRENT_STATE, NEXT_STATE:STATES;
BEGIN
    PROCESS (CLK)
    BEGIN
    IF CLK'EVENT AND CLK='1' THEN 
		CURRENT_STATE<=NEXT_STATE; 
		IF CURRENT_STATE=ST6 AND BUCKIN='0' THEN
		RESULT<='1';
		ELSE 
		RESULT<='0';
		END IF;
	 END IF;
    END PROCESS;
    PROCESS (BUCKIN)
    BEGIN
        CASE CURRENT_STATE IS
            WHEN ST0 => IF BUCKIN = '1' THEN NEXT_STATE <= ST1; ELSE NEXT_STATE <= ST0; END IF;
            WHEN ST1 => IF BUCKIN = '1' THEN NEXT_STATE <= ST2; ELSE NEXT_STATE <= ST0; END IF;
            WHEN ST2 => IF BUCKIN = '1' THEN NEXT_STATE <= ST3; ELSE NEXT_STATE <= ST0; END IF;
            WHEN ST3 => IF BUCKIN = '0' THEN NEXT_STATE <= ST4; ELSE NEXT_STATE <= ST0; END IF;
            WHEN ST4 => IF BUCKIN = '0' THEN NEXT_STATE <= ST5; ELSE NEXT_STATE <= ST0; END IF;
            WHEN ST5 => IF BUCKIN = '1' THEN NEXT_STATE <= ST6; ELSE NEXT_STATE <= ST0; END IF;
            WHEN ST6 => IF BUCKIN = '0' THEN NEXT_STATE <= ST0; ELSE NEXT_STATE <= ST0; END IF;
				WHEN OTHERS => NEXT_STATE <= ST0;
        END CASE;
END PROCESS;
END BHV;