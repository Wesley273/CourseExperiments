CIRCUIT EXP2_3
VX 0 3 0
R1 1 2 RMOD 10
C1 1 0 CMOD 5UF IC=10V
L1 1 0 LMOD 5UH
W1 3 2 VX SMOD
.MODEL RMOD RES(R=1 TCE=3)
.MODEL LMOD IND(L=1 IL1=0.1 IL2=0.01 TC1=0.01 TC2=0.002)
.MODEL CMOD CAP(C=1 VC1=0.1 VC2=0.03 TC1=0.01 TC2=0.002)
.MODEL SMOD ISWITCH (RON=0.01 ROFF=10E+6 ION=1MA IOFF=0.1MA) 
.TRAN 2US 200US UIC
.TEMP 60
.PROBE
.PRINT TRAN I(VX)
.END