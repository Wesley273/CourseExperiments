CIRCUIT EXP5_3
VAB 2 0 DC 2V
R1 1 2 RMOD 1
R2 3 2 RMOD 1
R3 3 4 RMOD 1
R4 3 0 RMOD 1
R5 2 6 RMOD 1
R6 1 5 RMOD 1
R7 5 8 RMOD 1
R8 0 8 RMOD 1
R9 6 0 RMOD 1
R10 4 8 RMOD 1
R11 5 6 RMOD 1
R12 4 1 RMOD 1
.MODEL RMOD RES(R=1)
.DC VAB 0V 10V 1V 
.PROBE
.END