CIRCUIT EXP5_5
IS 0 1 AC 1A
R1 1 0 1K
R2 1 2 1K
C1 1 0 1UF
C2 2 0 1UF
.AC LIN 100000 1MHZ 200KHZ
.PROBE
.END