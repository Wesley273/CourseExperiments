CIRCUIT EXP4_3
VI 1 0 SIN(0V 1V 1MEGHZ)
RI 1 0 RMOD 1MEG
R1 2 0 RMOD 1G
R2 3 4 RMOD 1K
RO 4 0 RMOD 1G
E1 3 0 VALUE={2*V(1)*V(2)}
G1 2 0 VALUE={1-V(1)*V(1)}
G2 0 2 VALUE={V(2)*V(2)}
.MODEL RMOD RES(R=1 TCE=0)
.TRAN 10N 4U 0 1N
.PROBE
.END