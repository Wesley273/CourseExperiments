CIRCUIT EXAM_6
.SUBCKT QNPN 6 7 5
V1 1 7 DC 0V
RB 1 2 100
RPI 2 3 1K
RU 2 4 1MEG
RE 3 5 1
RO 4 3 100K
RC 4 6 10
CU 2 4 1PF
CPI 2 3 2PF
CCS 6 0 2PF
F1 3 4 V1 20
.ENDS QNPN
VIN 1 0 AC 10MV 0DEG
VC 0 7 DC 15V
RS 1 2 500
R1 3 7 47K
R2 3 0 5K
RC 4 7 10K
RE 5 0 2K
RL 6 0 20K
C1 2 3 1UF
CE 5 0 10UF
C2 4 6 1UF
X1 4 3 5 QNPN
.AC LIN 100000 1HZ 20KHZ
.PROBE
.END
