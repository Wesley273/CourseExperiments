LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY TRAFFIC_vhd_tst IS
END TRAFFIC_vhd_tst;
ARCHITECTURE TRAFFIC_arch OF TRAFFIC_vhd_tst IS
	SIGNAL CLK1 : STD_LOGIC;
	SIGNAL GF1 : STD_LOGIC;
	SIGNAL GM1 : STD_LOGIC;
	SIGNAL RF1 : STD_LOGIC;
	SIGNAL RM1 : STD_LOGIC;
	SIGNAL RST1 : STD_LOGIC;
	SIGNAL YF1 : STD_LOGIC;
	SIGNAL YM1 : STD_LOGIC;
	COMPONENT TRAFFIC
		PORT (
			CLK : IN STD_LOGIC;
			GF : OUT STD_LOGIC;
			GM : OUT STD_LOGIC;
			RF : OUT STD_LOGIC;
			RM : OUT STD_LOGIC;
			RST : IN STD_LOGIC;
			YF : OUT STD_LOGIC;
			YM : OUT STD_LOGIC
		);
	END COMPONENT;
	CONSTANT CLK_P : TIME := 500 MS;
BEGIN
	i1 : TRAFFIC
	PORT MAP(
		CLK => CLK1,
		GF => GF1,
		GM => GM1,
		RF => RF1,
		RM => RM1,
		RST => RST1,
		YF => YF1,
		YM => YM1
	);

	PROCESS BEGIN
		CLK1 <= '0';
		WAIT FOR CLK_P;
		CLK1 <= '1';
		WAIT FOR CLK_P;
	END PROCESS;
	RST1 <= '1', '0' AFTER 3000 MS;
END TRAFFIC_arch;