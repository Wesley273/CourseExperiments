LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY ELEVATOR_vhd_tst IS
END ELEVATOR_vhd_tst;
ARCHITECTURE ELEVATOR_arch OF ELEVATOR_vhd_tst IS
	SIGNAL CLK1 : STD_LOGIC;
	SIGNAL DOOR_LIGHT1 : STD_LOGIC;
	SIGNAL DOWN1 : STD_LOGIC_VECTOR(10 DOWNTO 1);
	SIGNAL INSIDE1 : STD_LOGIC_VECTOR(10 DOWNTO 1);
	SIGNAL POSITION1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL RST1 : STD_LOGIC;
	SIGNAL UP1 : STD_LOGIC_VECTOR(10 DOWNTO 1);
	COMPONENT ELEVATOR
		PORT (
			CLK : IN STD_LOGIC;
			DOOR_LIGHT : OUT STD_LOGIC;
			DOWN : IN STD_LOGIC_VECTOR(10 DOWNTO 1);
			INSIDE : IN STD_LOGIC_VECTOR(10 DOWNTO 1);
			POSITION : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			RST : IN STD_LOGIC;
			UP : IN STD_LOGIC_VECTOR(10 DOWNTO 1)
		);
	END COMPONENT;
	CONSTANT CLK_P : TIME := 500 MS;
BEGIN
	i1 : ELEVATOR
	PORT MAP(
		CLK => CLK1,
		DOOR_LIGHT => DOOR_LIGHT1,
		DOWN => DOWN1,
		INSIDE => INSIDE1,
		POSITION => POSITION1,
		RST => RST1,
		UP => UP1
	);
	PROCESS BEGIN
		CLK1 <= '0';
		WAIT FOR CLK_P;
		CLK1 <= '1';
		WAIT FOR CLK_P;
	END PROCESS;
	RST1 <= '1', '0' AFTER 200 MS;
	INSIDE1 <= "0000000000", "0000010000" AFTER 5000 MS, "0000000000" AFTER 11000 MS, "0010000000" AFTER 19000 MS, "0000100000" AFTER 32000 MS, "0000000000" AFTER 50000 MS;
	UP1 <= "0001000100", "0000000000" AFTER 35000 MS;
	DOWN1 <= "0100000000", "0000000000" AFTER 35000 MS;
END ELEVATOR_arch;