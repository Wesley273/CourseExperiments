CIRCUIT EXP8_3
.LIB C:\Users\Wesley\Documents\Git\ElectronicDesign\PSpice\EXP8\my_lib.lib
.SUBCKT COMPARER 3 2 4 8 7
VB 10 0 DC 1.85V
VE 0 12 DC 1.85V
IEE 5 4 DC 0.4MA
IOS 0 14 DC 9.25MA
IO 7 4 DC 2.5MA
GA 9 0 VALUE={(2.3E-4)*(V(15)-V(6))}
GB 11 0 VALUE={(7.8E-5)*(V(15)-V(6))}
GC 14 0 VALUE={(5E-3)*V(9)}
RC1 8 6 10K
RC2 15 8 10K
RPC 8 0 2.5K
RPE 4 0 3.5K
RA 9 0 100K
RB 11 0 300K
RO 14 0 200
C1 9 0 0.56PF
Q1 6 2 5 QN1
Q2 15 3 5 QN1
D1 6 15 DN1
D2 15 6 DN2
D3 9 10 DN3
D4 12 9 DN3
D5 9 11 DN3
D6 14 7 DN3
.ENDS
VREF1 1 0 DC 4V
VREF2 3 0 DC -4V
VIN 2 0 DC 1V
VCC 11 0 DC 12V
VEE 10 0 DC -6V
R1 1 4 10K
R2 10 7 2K
R3 2 5 5K
R4 3 6 10K
R5 10 8 2K
R6 9 0 10K
D1 7 9 DN4
D2 8 9 DN4
X1 4 5 10 11 7 COMPARER
X2 5 6 10 11 8 COMPARER
.DC VIN -10V 10V 0.01V
.PROBE
.END
