CIRCUIT EXP4_9
VS 3 0 PWL(0 1V 1NS 1V 1.001US 0V)
VI 1 0 PWL(0 0V 100US 1V 200US 1V 210US 2V 300US 2V 310US 3V 400US 3V)
VBH 5 0 DC 1V
VBL 0 6 DC 1V
RI 1 0 RMOD 1E+6
R1 2 0 RMOD 1T
R2 4 0 RMOD 1K
CT 3 2 1NF
C2 4 0 100PF
D1 4 5 DMOD
D2 6 4 DMOD
G1 0 2 POLY(2) 4 0 1 0 0 -2E-4 0 0 -1E-4
G2 0 4 POLY(2) 2 0 4 0 0 1 1
.MODEL RMOD RES(R=1 TCE=0)
.MODEL DMOD D N=0.01
.OPTIONS ITL5=0
.TRAN 1US 400U
.PROBE
.END