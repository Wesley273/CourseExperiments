LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY HADDER1 IS
        PORT (
                A, B : IN STD_LOGIC;
                CO : OUT STD_LOGIC;
                SO : OUT STD_LOGIC
        );
END HADDER1;
ARCHITECTURE ONE OF HADDER1 IS
BEGIN
        SO <= A XOR B;
        CO <= A AND B;
END ONE;