CIRCUIT EXP8_1
VI 1 0 DC 1V
VZ 0 4 DC 12V
R1 1 2 0.001
R2 2 3 RMOD 0.1
D1 2 0 DMOD2
D2 4 3 DMOD1
.MODEL RMOD RES(R=1)
.MODEL DMOD1 D N=0.001
.MODEL DMOD2 D
.DC VI -13V -10V 0.01V
.STEP RES RMOD(R) LIST 1 10 100
*.STEP VZ LIST 6V 8V 10V
.PROBE
.END
