LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY GATE_OR IS
       PORT (
              A, B : IN STD_LOGIC;
              C : OUT STD_LOGIC
       );
END GATE_OR;
ARCHITECTURE ONE OF GATE_OR IS
BEGIN
       C <= A OR B;
END ONE;