CIRCUIT EXP2_2
R1 2 3 RMOD 10
R2 1 4 RMOD 10K
R3 0 5 RMOD 5K
C1 4 0 CMOD 100UF
C2 0 5 CMOD 10UF
L1 3 0 1H
L2 0 1 15MH
L3 5 0 15MH
KALL L1 L2 L3 0.9999
V1 2 0 SIN(0 220 50)
.MODEL RMOD RES (R=2 TC1=0.2 TC2=2.5)
.MODEL CMOD CAP (C=2 VC1=0.05 VC2=0.015 TC1=0.02 TC2=0.006)
.TRAN 0.1M 60M 0 0.01M
.TEMP 50
.PRINT TRAN V(5)
.PROBE
.END