LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ADDER4 IS
     PORT (
          CIN : IN STD_LOGIC;
          A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
          B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
          SUM : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
          COUT : OUT STD_LOGIC);
END ENTITY ADDER4;

ARCHITECTURE ART OF ADDER4 IS
     SIGNAL S5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
     SIGNAL A5, B5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
     A5 <= '0' & A;
     B5 <= '0' & B;
     S5 <= A5 + B5 + CIN;
     SUM <= S5(3 DOWNTO 0);
     COUT <= S5(4);
END ARCHITECTURE ART;