LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY COMPARER4 IS
	PORT (
		A3 : IN STD_LOGIC;
		A2 : IN STD_LOGIC;
		A1 : IN STD_LOGIC;
		A0 : IN STD_LOGIC;
		B3 : IN STD_LOGIC;
		B2 : IN STD_LOGIC;
		B1 : IN STD_LOGIC;
		B0 : IN STD_LOGIC;
		G : OUT STD_LOGIC;
		M : OUT STD_LOGIC;
		L : OUT STD_LOGIC
	);
END ENTITY COMPARER4;
ARCHITECTURE BHV OF COMPARER4 IS
	SIGNAL INDATAA : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL INDATAB : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	INDATAA <= A3 & A2 & A1 & A0;
	INDATAB <= B3 & B2 & B1 & B0;
	P1 : PROCESS (A3, A2, A1, A0, B3, B2, B1, B0)
	BEGIN
		IF (INDATAA > INDATAB) THEN
			G <= '1';
			M <= '0';
			L <= '0';
		ELSIF (INDATAA = INDATAB) THEN
			M <= '1';
			L <= '0';
			G <= '0';
		ELSIF (INDATAA < INDATAB) THEN
			L <= '1';
			G <= '0';
			M <= '0';
		END IF;
	END PROCESS P1;
END BHV;