CIRCUIT EXP3_1
*VI 3 0 EXP (0.5 10 2US 2US 10US 2US)
*VI 3 0 PULSE(0.2V 5V 1US 3US 1US 10US 16US)
VI 3 0 PWL(0 0.1V 3US 0.1V 5US 1V 8US 3V 9US 5V 13US 1V 15US 0.1V)
V1 6 0 DC 12V
V2 0 9 DC 12V
R1 0 4 RMOD 5.6K
R7 11 6 RMOD 1K
R8 2 9 RMOD 1K
C1 1 4 CMOD 100UF
C2 4 0 CMOD 100PF
L1 4 0 LMOD 10UH
D1 11 3 DMOD
D2 3 2 DMOD
Q1 6 11 1 QNPN
Q2 9 2 1 QPNP
.MODEL RMOD RES(R=1 TCE=0)
.MODEL LMOD IND(L=1 IL1=0 IL2=0 TC1=0 TC2=0)
.MODEL CMOD CAP(C=1 VC1=0 VC2=0 TC1=0 TC2=0)
.MODEL DMOD D IS=2E-13 RS=5 N=2
.MODEL QNPN NPN(IS=5E-10 BF=250 RB=50 VAF=100)
.MODEL QPNP PNP(IS=5E-10 BF=250 RB=50 VAF=100)
.TRAN 1US 20US
.PROBE
.END