CIRCUIT EXAM_3
.LIB C:\Users\Wesley\Documents\Git\ElectronicDesign\PSpice\EXAM\eval.lib
VI1 1 0 DC {VE}
VI2 2 0 DC {6-VE}
VCC 5 0 DC 15V
VSS 6 0 DC -15V
R1 2 3 10K
R2 3 0 5K
R3 3 4 10K
X1 1 3 5 6 4 uA741
.PARAM VE=(TEMP-5)/2
.DC PARAM VE 0V 4V 0.1V
.PROBE
.END