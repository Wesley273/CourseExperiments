CIRCUIT EXP4_5
VCC 1 0 DC 5V
RR 1 2 RMOD 1K
R0 3 0 RMOD 1K
R1 4 0 RMOD 2K
R2 5 0 RMOD 1K
R3 6 0 RMOD 0.5K
Q0 1 2 3 QNPN
Q1 1 2 4 QNPN
Q2 1 2 5 QNPN
Q3 1 2 6 QNPN
.MODEL RMOD RES(R=1 TCE=0)
.MODEL QNPN NPN
.TRAN 10U 4M
.PROBE
.END