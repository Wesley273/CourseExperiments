CIRCUIT EXAM_4
V1 1 0 DC 1V
R1 3 1 3
R2 1 0 1
R3 3 0 1
R4 3 4 3
R5 0 4 1
R6 1 4 3
.TRAN 0 1000US
.PROBE
.END