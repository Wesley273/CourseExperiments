CIRCUIT EXP5_1
V1 8 0 DC 0V AC 1V 30DEG SFFM (0.2V 0.1V 10KHZ 5 1KHZ)
VC 3 0 DC 12V
R1 1 2 10K
R2 1 3 RMOD 1K
RB2 2 0 20K
RC1 3 4 3K
RE1 5 0 2K
RL1 6 0 3K
C1 8 2 10UF
C2 4 6 10UF IC=0.1V
CE1 5 0 47UF
Q1 4 2 5 QNPN
.MODEL RMOD RES(R=57)
.MODEL QNPN NPN(IS=2.5E-15A BF=250 RB=300 VAF=100 Cjc=3.638pF Cje=4.493pF)

*******DC Analysis*******
*.DC RES RMOD(R) 1 100 1
*************************

*******AC Analysis*******
*.AC DEC 10 1MEGHZ 10MEGHZ
*************************

****Transient Analysis****
*.TRAN 1US 100US UIC
**************************

.SENS V(4)
.PROBE
.END