CIRCUIT EXP3_6
VA 1 0 PWL(0 0V 1NS 0V 2NS 3.6V 20US 3.6V 20.001US 0V)
VB 2 0 DC 3.6V
VC 3 0 DC 3.6V
VCC 11 0 DC 5V
R1 4 11 RMOD 2.8K
R2 6 11 RMOD 750
R3 7 8 RMOD 300
R4 12 11 RMOD 75
R5 9 0 RMOD 3K
R6 7 10 RMOD 200
R11 11 14 RMOD 2.8K
D1 15 16 DMOD
D2 16 0 DMOD
Q1A 5 4 1 QNPN
Q1B 5 4 2 QNPN
Q1C 5 4 3 QNPN
Q2 6 5 7 QNPN
Q3 12 6 9 QNPN
Q4 12 9 13 QNPN
Q5 13 7 0 QNPN
Q6 10 8 0 QNPN
Q11 15 14 13 QNPN
.MODEL RMOD RES(R=1 TCE=0)
.MODEL DMOD D(IS=5E-14 RS=5 TT=0.1NS)
.MODEL QNPN NPN(IS=5E-14 BF=60 RB=60 RC=20 VAF=60 CJC=4P TF=0.1NS TR=10NS)
.TRAN 0.1US 45US
.PROBE
.END