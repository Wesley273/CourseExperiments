CIRCUIT EXP4_2
V1 1 0 DC 12V
VX 6 4 DC 0V
I1 4 2 DC 1A
R1 1 2 RMOD 2
R2 3 0 RMOD 2
R3 2 6 RMOD 2
R4 4 0 RMOD 2
R5 4 5 RMOD 2
H1 2 3 VX 0.2
G1 5 0 VALUE={0.1*V(3)}
.MODEL RMOD RES(R=1 TCE=0)
.TRAN 10N 4U 0 1N
.PROBE
.OP
.END