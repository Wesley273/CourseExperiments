CIRCUIT EXP5_8
V1 1 0 PWL(0S 2V 1S 2V 1.000001S 0V 2S 0V)
V2 2 0 PWL(0S 0V 1S 0V 1.000001S 2V 2S 2V)
VS 3 0 DC 10V
R1 6 4 10
R2 4 5 10
R3 5 0 10
R4 1 0 1E9
R5 2 0 1E9
L1 5 0 1H
S1 3 6 1 0 SMOD
S2 4 0 2 0 SMOD
.MODEL SMOD VSWITCH (RON=0.01 ROFF=1E+9 VON=1V VOFF=0V) 
.TRAN 1S 2S 
.PROBE
.END