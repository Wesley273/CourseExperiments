LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CNT10_DECODE IS
    PORT (
        CLK, RST, EN, LOAD : IN STD_LOGIC;
        DATA : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        DOUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        COUT : OUT STD_LOGIC;
        SG_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END CNT10_DECODE;
ARCHITECTURE BHV OF CNT10_DECODE IS
    COMPONENT FDIVIDER IS
        PORT (
            CLK : IN STD_LOGIC; --50MHz
            CP2 : BUFFER STD_LOGIC := '0';
            CP1 : BUFFER STD_LOGIC := '0');
    END COMPONENT FDIVIDER;
    COMPONENT CNT10 IS
        PORT (
            CLK, RST, EN, LOAD : IN STD_LOGIC;
            DATA : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            DOUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            COUT : OUT STD_LOGIC);
    END COMPONENT CNT10;
    COMPONENT DECODER7 IS
        PORT (
            BIN_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            SG_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    END COMPONENT DECODER7;
    SIGNAL CLKIN : STD_LOGIC;
    SIGNAL TOSG : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
BEGIN
    GETCLK : FDIVIDER PORT MAP(CLK => CLK, CP1 => CLKIN);
    COUNTER : CNT10 PORT MAP(CLK => CLKIN, RST => RST, EN => EN, LOAD => LOAD, DATA => DATA, DOUT => TOSG(3 DOWNTO 0), COUT => TOSG(4));
    DECODER_HIGH : DECODER7 PORT MAP(BIN_IN => TOSG(7 DOWNTO 4), SG_OUT => SG_OUT(15 DOWNTO 8));
    DECODER_LOW : DECODER7 PORT MAP(BIN_IN => TOSG(3 DOWNTO 0), SG_OUT => SG_OUT(7 DOWNTO 0));
    DOUT <= TOSG(3 DOWNTO 0);
    COUT <= TOSG(4);
END BHV;