R2 0 2 33K
R3 4 0 5.6K
L1 4 0 LMOD 10UH IC=1A
C1 2 0 CMOD 100UF IC=1V
C2 3 4 CMOD 100UF
C3 0 4 CMOD 100PF
S1 2 3 2 0 SMOD
.MODEL LMOD IND(L=1 IL1=0.3 IL2=0.005 TC1=0 TC2=0)
.MODEL CMOD CAP(C=1 VC1=0.05 VC2=0.01 TC1=0 TC2=0)
.MODEL SMOD VSWITCH(RON=5E-3 ROFF=1E+7 VON=0.7V VOFF=0)

.TRAN  2US 100US  UIC
.PROBE
.PRINT TRAN I(R3)
.END
