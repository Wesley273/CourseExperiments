CIRCUIT EXP6_2
.LIB C:\Users\Wesley\Documents\PSpice\EXP6\eval.lib

.SUBCKT INVERTER 1 2 3 4
* NODES: VDD,VIN,VOUT,VSS 
M1 3 2 1 1 IRF9140
M2 3 2 4 4 IRF150
C1 3 4 1UF
.ENDS INVERTER

VDD 4 0 DC 5V
X1 4 1 2 0 INVERTER
X2 4 2 3 0 INVERTER
X3 4 3 1 0 INVERTER
.TRAN 10US 30US
.IC V(1)=0
.PROBE
.END
