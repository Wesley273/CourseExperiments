CIRCUIT EXP7_2
.SUBCKT AMPLIFIRE 1 2 7 9 8
R1 6 9 140K
C1 8 4 CMOD 1.6PF
M1 3 1 5 5 MOD1 W=30U L=20U AD=200P AS=200P
M2 4 2 5 5 MOD1 W=30U L=20U AD=200P AS=200P
M3 3 3 9 9 MOD2 W=50U L=12U AD=300P AS=300P
M4 4 3 9 9 MOD2 W=50U L=12U AD=300P AS=300P
M5 5 6 7 7 MOD1 W=80U L=20U AD=400P AS=400P
M6 6 6 7 7 MOD1 W=40U L=20U AD=300P AS=300P
M7 8 4 9 9 MOD2 W=198U L=12U AD=500P AS=500P
M8 8 6 7 7 MOD1 W=158U L=20U AD=400P AS=400P
.MODEL MOD1 PMOS(
+LEVEL=2 VTO=-1.0 LAMBDA=0.005 
+PB=0.98 CGSO=2.88E-9 CGDO=2.88E-9 CGBO=1.38E-9 
+RSH=100 CJ=2.2E-4 MJ=0.5 JS=0.01 TOX=8E-8 
+NSUB=5E15 TPG=-1 XJ=1E-6 LD=0.6U UO=200 
+UCRIT=6E4 UEXP=0.15 UTRA=0.3 
+VMAX=5E4 NEFF=3 XQC=0.4 DELTA=8
)
.MODEL MOD2 NMOS(
+LEVEL=2 VTO=1.0 LAMBDA=0.005 
+PB=0.98 CGSO=2.88E-9 CGDO=2.88E-9 CGBO=1.38E-9 
+RSH=20 CJ=4.3E-4 MJ=0.5 JS=0.01 TOX=8E-8 
+NSUB=2E16 TPG=1 XJ=1E-6 LD=0.6U UO=600 
+UCRIT=6E4 UEXP=0.2 UTRA=0.3 
+VMAX=5E4 NEFF=3 XQC=0.4 DELTA=8
)
.MODEL CMOD CAP(C=1)
.ENDS

V1 6 0 SIN(0V 100MV 5KHZ)
V2 7 0 PULSE(-1V 1V 0 1NS 1NS 0.5MS 1MS)
VDD 4 0 DC 7.5V
VSS 5 0 DC -7.5V
R1 7 1 15K
R2 6 1 15K
R3 2 3 30K
R4 2 0 10K
X1 2 1 4 5 3 AMPLIFIRE
.TRAN 1MS 2MS
.PROBE
.END
