CIRCUIT EXP4_7
V1 1 0 SIN(0V 1V 1KHZ)
V2 2 0 SIN(0V 1V 1KHZ)
V3 3 0 SIN(0V 1V 1KHZ)
R1 1 0 RMOD 1
R2 2 0 RMOD 2
R3 3 0 RMOD 5
RO 5 4 RMOD 1K
RL 5 0 RMOD 1G
*H1 4 0 POLY(3) V1 V2 V3 0 0 0 1 1 0 0 1 0 1
E1 4 0 VALUE={I(V3)+I(V1)*I(V1)+I(V2)*I(V2)+I(V3)*I(V3)}
.MODEL RMOD RES(R=1 TCE=0)
.TRAN 20U 2M
.PROBE
.END