CIRCUIT EXP4_1
V1 1 0 SIN(0V 1V 5KHZ)
V2 2 0 SIN(1V 0.9V 1KHZ)
R1 1 0 RMOD 1G
R2 2 0 RMOD 1G
RL 3 0 RMOD 1MEG
E1 3 0 POLY(2) 1 0 2 0 0 0 0 0 1
.MODEL RMOD RES(R=1 TCE=0)
.TRAN 1U 0.8M
.PROBE
.OP
.END