CIRCUIT EXAM_5
I1 0 7 DC 1A
I2 6 3 DC 1A
I3 0 3 DC 3A
I4 9 2 DC 3A
I5 2 3 DC 2A
V1 8 9 DC 10V
V2 4 3 DC 10V
V3 2 1 DC 6V
V4 10 2 DC 4V
R1 6 8 4
R2 7 4 2
R3 1 0 3
R4 3 10 1
R5 3 6 1G
R6 2 9 1G
.TRAN 0 100US
.SENS I(V4)
.PROBE
.END