CIRCUIT EXP4_4
VI 2 0 SIN(0V 10V 1KHZ)
VS1 1 0 DC 0V
VS2 3 0 DC 0V
F1 0 2 VS2 4
F2 0 4 VS1 0.25
R1 2 1 RMOD 2K
R2 3 4 RMOD 8K
RL 4 0 RMOD 8K
.MODEL RMOD RES(R=1 TCE=0)
.TRAN 10U 4M
.PROBE
.END