CIRCUIT EXP7_1
VDD 7 0 DC 7.5V
VSS 9 0 DC -7.5V
VI1 1 0 DC 0V
VI2 2 0 AC 1V
R1 6 9 140K
C1 8 4 CMOD 1.6PF
M1 3 1 5 5 MOD1 W=30U L=20U AD=200P AS=200P
M2 4 2 5 5 MOD1 W=30U L=20U AD=200P AS=200P
M3 3 3 9 9 MOD2 W=50U L=12U AD=300P AS=300P
M4 4 3 9 9 MOD2 W=50U L=12U AD=300P AS=300P
M5 5 6 7 7 MOD1 W=80U L=20U AD=400P AS=400P
M6 6 6 7 7 MOD1 W=40U L=20U AD=300P AS=300P
M7 8 4 9 9 MOD2 W=198U L=12U AD=500P AS=500P
M8 8 6 7 7 MOD1 W=158U L=20U AD=400P AS=400P
.MODEL MOD1 PMOS(
+LEVEL=2 VTO=-1.0 LAMBDA=0.005 
+PB=0.98 CGSO=2.88E-9 CGDO=2.88E-9 CGBO=1.38E-9 
+RSH=100 CJ=2.2E-4 MJ=0.5 JS=0.01 TOX=8E-8 
+NSUB=5E15 TPG=-1 XJ=1E-6 LD=0.6U UO=200 
+UCRIT=6E4 UEXP=0.15 UTRA=0.3 
+VMAX=5E4 NEFF=3 XQC=0.4 DELTA=8
)
.MODEL MOD2 NMOS(
+LEVEL=2 VTO=1.0 LAMBDA=0.005 
+PB=0.98 CGSO=2.88E-9 CGDO=2.88E-9 CGBO=1.38E-9 
+RSH=20 CJ=4.3E-4 MJ=0.5 JS=0.01 TOX=8E-8 
+NSUB=2E16 TPG=1 XJ=1E-6 LD=0.6U UO=600 
+UCRIT=6E4 UEXP=0.2 UTRA=0.3 
+VMAX=5E4 NEFF=3 XQC=0.4 DELTA=8
)
.MODEL CMOD CAP(C=1)
.STEP CAP CMOD(C) LIST 1.6 5 10
.AC DEC 1HZ 100 10MEGHZ 
.TEMP 27
.PROBE
.END