LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY WORK;
ENTITY MUX41 IS
	PORT (
		S0 : IN STD_LOGIC;
		D2 : IN STD_LOGIC;
		INH : IN STD_LOGIC;
		D0 : IN STD_LOGIC;
		D1 : IN STD_LOGIC;
		D3 : IN STD_LOGIC;
		S1 : IN STD_LOGIC;
		Q : OUT STD_LOGIC
	);
END MUX41;

ARCHITECTURE BDF_TYPE OF MUX41 IS

	SIGNAL SYNTHESIZED_WIRE_18 : STD_LOGIC;
	SIGNAL SYNTHESIZED_WIRE_19 : STD_LOGIC;
	SIGNAL SYNTHESIZED_WIRE_20 : STD_LOGIC;
	SIGNAL SYNTHESIZED_WIRE_21 : STD_LOGIC;
	SIGNAL SYNTHESIZED_WIRE_22 : STD_LOGIC;
	SIGNAL SYNTHESIZED_WIRE_13 : STD_LOGIC;
	SIGNAL SYNTHESIZED_WIRE_14 : STD_LOGIC;
	SIGNAL SYNTHESIZED_WIRE_15 : STD_LOGIC;
	SIGNAL SYNTHESIZED_WIRE_16 : STD_LOGIC;

BEGIN
	SYNTHESIZED_WIRE_18 <= NOT(S0);
	SYNTHESIZED_WIRE_21 <= NOT(SYNTHESIZED_WIRE_18);
	SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_18 AND D0;
	SYNTHESIZED_WIRE_14 <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_21 AND D1;
	SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_22 AND SYNTHESIZED_WIRE_18 AND D2;
	SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_22 AND SYNTHESIZED_WIRE_21 AND D3;
	Q <= SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15 OR SYNTHESIZED_WIRE_16;
	SYNTHESIZED_WIRE_19 <= NOT(INH);
	SYNTHESIZED_WIRE_20 <= NOT(S1);
	SYNTHESIZED_WIRE_22 <= NOT(SYNTHESIZED_WIRE_20);
END;