CIRCUIT EXAM_2
V1 1 0 PULSE(1V 5V 1MS 2MS 2MS 3MS 10MS)
R1 1 2 RMOD 4
C1 1 2 CMOD 100UF
L1 2 3 LMOD 0.02H
C2 3 4 CMOD 50UF
R2 4 0 RMOD 3
.MODEL RMOD RES(R=1 TC1=0.002 TC2=0.005)
.MODEL CMOD CAP(C=1 TC1=0.01 TC2=0.002)
.MODEL LMOD IND(L=1 TC1=0.02 TC2=0.003)
.TEMP 10 27 32
.TRAN 5MS 15MS
.PROBE
.END