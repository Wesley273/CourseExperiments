CIRCUIT EXP6_1
V1 7 0 SIN(0V 100MV 1KHZ)
VCC 9 0 DC 12V
VEE 10 0 DC -12V
R1 1 9 RMOD 10K
R2 2 9 RMOD 10K
R3 3 10 RMOD 10K
R4 5 9 RMOD 300K
R5 6 9 RMOD 300K
R6 7 5 RMOD 2K
R7 7 6 RMOD 2K
R8 8 0 RMOD 1G
R9 4 0 RMOD 1G
C1 1 8 CMOD 10UF
C2 4 2 CMOD 10UF
Q1 1 5 3 QNPN
Q2 2 6 3 QNPN
.MODEL RMOD RES(R=1 DEV=30% LOT=20%)
.MODEL CMOD CAP(C=1 DEV=20% LOT=10%)
.MODEL QNPN NPN(BF=200 DEV=20%)
.TRAN 10US 2MS
*******MC Analysis*******
*.MC 10 TRAN V(8,4) YMAX LIST OUTPUT ALL
*************************

*******WCASE Analysis*******
.WCASE TRAN V(8) YMAX DEVICES QNPN
****************************
.PROBE
.END
