CIRCUIT EXP7_6
V1 1 0 AC 1V 0DEG
R1 1 2 1
L1 2 3 1E-4H
C1 3 0 100UF
R2 3 0 1
.AC LIN 1000 1590HZ 1592HZ
.PROBE
.END