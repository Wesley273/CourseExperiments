LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ADDER16_B_vhd_tst IS
END ADDER16_B_vhd_tst;
ARCHITECTURE ADDER16_B_arch OF ADDER16_B_vhd_tst IS
	SIGNAL A1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL B1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL CIN1 : STD_LOGIC;
	SIGNAL COUT1 : STD_LOGIC;
	SIGNAL SUM1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
	COMPONENT ADDER16_B
		PORT (
			A : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			CIN : IN STD_LOGIC;
			COUT : OUT STD_LOGIC;
			SUM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
BEGIN
	i1 : ADDER16_B
	PORT MAP(
		A => A1,
		B => B1,
		CIN => CIN1,
		COUT => COUT1,
		SUM => SUM1
	);
	A1 <= "1100111100001111", "1000000011110000" AFTER 100 NS, "0111111100100111" AFTER 800 NS;
	B1 <= "1100111100001100", "1000110000001100" AFTER 100 NS, "0110011111111111" AFTER 800 NS;
	CIN1 <= '1', '0' AFTER 500 NS, '1' AFTER 800NS;
END ADDER16_B_arch;