CIRCUIT EXP5_6
VCC 5 0 DC 6V
RC1 5 2 3K
RB2 5 3 40K
RB1 5 1 40K
RC2 5 6 3K
C1 2 3 100PF
C2 1 6 100PF
Q1 2 1 0 QNPN
Q2 6 3 0 QNPN
.MODEL QNPN NPN(IS=2E-15A BF=80 RB=10 RC=5 TF=10NS CJC=1PF CJE=1PF)
.TRAN 20US 100US UIC
.IC V(1)=0V
.IC V(2)=6V
.PROBE
.END