CIRCUIT EXP3_3
VS 1 0 16V
IS 3 4 1A
R2 4 0 RMOD 3
R3 2 3 RMOD 4
R4 3 0 RMOD 20
R5 1 2 RMOD 8
RL 2 4 RMOD 3
.MODEL RMOD RES(R=1 TCE=0)
.DC VS 0 16 8
.PRINT DC I(RL)
.END