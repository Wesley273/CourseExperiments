CIRCUIT EXP5_4
VG 1 0 DC 2V
VD 2 0 DC 2V
M1 2 1 0 0 MNMOS
.MODEL RMOD RES(R=1)
.MODEL MNMOS NMOS(IS=1E-32 VTO=1 LAMBDA=0.0457468 KP=179.181 CGSO=5.51447E-05 CGDO=1E-11)
.DC VG 2V 6V 1V 
.PROBE
.END