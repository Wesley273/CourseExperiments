CIRCUIT EXP7_4
VS 2 1 SIN(0V {VA(X1)} 1KHZ)
VBB 1 0 DC 0.7V
VCC 4 0 DC 12V
RC 4 3 2K
Q1 3 2 0 QNPN
.MODEL QNPN NPN(IS=2E-15  BF=200  RB=60)
.FUNC VA(X) {(2*X-5MV)}
.PARAM X1=5MV
.TRAN 0MS 0.3MS 0.01MS
.STEP PARAM X1 LIST 5MV 7.5MV 10MV 12.5MV 15MV
.PROBE
.END