CIRCUIT EXP3_4
V1 1 7 AC 100MV 0DEG
V2 8 0 DC 15V
R1 4 8 RMOD 15K
R2 3 8 RMOD 1.4E+6
R3 3 0 RMOD 1E+6
R4 1 2 RMOD 250
R5 5 9 RMOD 100
R6 9 0 RMOD 15K
R7 6 7 RMOD 15K
R8 7 0 RMOD 5K
R9 6 0 RMOD 10K
C1 2 3 CMOD 1UF
C2 4 6 CMOD 0.1UF
C3 9 0 CMOD 20UF
M1 4 3 5 5 MNMOS
.MODEL RMOD RES(R=1 TCE=0)
.MODEL LMOD IND(L=1 IL1=0 IL2=0 TC1=0 TC2=0)
.MODEL CMOD CAP(C=1 VC1=0 VC2=0 TC1=0 TC2=0)
.MODEL MNMOS NMOS (VTO=1 KP=6.5E-3 CBD=5PF CBS=2PF RD=5 RS=2 RB=0 RG=0 RDS=1MEG CGSO=1PF CGDO=1PF CGBO=1PF)
.AC DEC 10 10HZ 100MEGHZ
.PRINT AC VM(7)
.OP
.PROBE
.END